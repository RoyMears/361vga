`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Roy Mears, Jonathan Zavala, Luis Arevalo
// 
// Create Date: 10/9/2023 5:28:33 AM
// Design Name: 
// Module Name: pongGraphicalAnimation
// Project Name: CECS361FinalProjectPong
// Target Devices: nexys a7 100t
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module pongGraphicalAnimation(

    );
    
    // can do majority of pixel generation here, or outsourse for objects
endmodule
